module fix_float_multiplier_tb (
    ports
);
    
endmodule 