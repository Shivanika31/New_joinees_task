module tb;
gggg
endmodule